module top_d1p1_tb
  
endmodule

module top_t1p1

endmodule
